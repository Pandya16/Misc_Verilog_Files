`timescale 1ns / 1ps
module bus16bit(o, d3, d2, d1, d0, s);
output [15:0] o;
input [15:0] d3;
input [15:0] d2;
input [15:0] d1;
input [15:0] d0;
input [1:0] s;
mux_4to1 x0(o[0],d0[0],d1[0],d2[0],d3[0],s[1:0]);
mux_4to1 x1(o[1],d0[1],d1[1],d2[1],d3[1],s[1:0]);
mux_4to1 x2(o[2],d0[2],d1[2],d2[2],d3[2],s[1:0]);
mux_4to1 x3(o[3],d0[3],d1[3],d2[3],d3[3],s[1:0]);
mux_4to1 x4(o[4],d0[4],d1[4],d2[4],d3[4],s[1:0]);
mux_4to1 x5(o[5],d0[5],d1[5],d2[5],d3[5],s[1:0]);
mux_4to1 x6(o[6],d0[6],d1[6],d2[6],d3[6],s[1:0]);
mux_4to1 x7(o[7],d0[7],d1[7],d2[7],d3[7],s[1:0]);
mux_4to1 x8(o[8],d0[8],d1[8],d2[8],d3[8],s[1:0]);
mux_4to1 x9(o[9],d0[9],d1[9],d2[9],d3[9],s[1:0]);
mux_4to1 x10(o[10],d0[10],d1[10],d2[10],d3[10],s[1:0]);
mux_4to1 x11(o[11],d0[11],d1[11],d2[11],d3[11],s[1:0]);
mux_4to1 x12(o[12],d0[12],d1[12],d2[12],d3[12],s[1:0]);
mux_4to1 x13(o[13],d0[13],d1[13],d2[13],d3[13],s[1:0]);
mux_4to1 x14(o[14],d0[14],d1[14],d2[14],d3[14],s[1:0]);
mux_4to1 x15(o[15],d0[15],d1[15],d2[15],d3[15],s[1:0]);
endmodule
