`timescale 1ns / 1ps
module mux_4to1(o, i1, i2, i3, i4, s);
output o;
input i1;
input i2;
input i3;
input i4;
input [1:0] s;
wire [5:0] m;

endmodule